package axi_pkg;
  import uvm_pkg::*;

  `include "uvm_macros.svh"
  `include "axi_include.svh"

endpackage
